`default_nettype none
`include "m_proc5.v"

module m_top();
  reg r_clk=0; initial #150 forever #50 r_clk = ~r_clk;
  reg [31:0] r_cc=1; always @(posedge r_clk) r_cc <= r_cc + 1;
  initial #1000000 begin $display("time out"); $finish; end
  m_proc5 m (r_clk);
  initial begin
    m.m3.mem[0]={12'd5,5'd0,3'h0,5'd1,7'h13};          //  addi x1,x0,5
    m.m3.mem[1]={7'd0,5'd1,5'd1,3'h0,5'd2,7'h33};      //  add  x2,x1,x1
    m.m3.mem[2]={12'd1,5'd1,3'h0,5'd1,7'h13};          //L:addi x1,x1,1
    m.m3.mem[3]={~7'd0,5'd2,5'd1,3'h1,5'b11101,7'h63}; //  bne  x1,x2,L
    m.m3.mem[4]={12'd9,5'd1,3'h0,5'd10,7'h13};         //  addi x10,x1,9
    m.m3.mem[5]=32'h00050f13;                          //  HALT
  end
  initial #99 forever #100 $display("CC%02d %h %d %d %d",
    r_cc, m.r_pc, m.w_r1, m.w_s2, m.w_rt);
endmodule
