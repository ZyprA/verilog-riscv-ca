module m_mux(w_in1, w_in2, w_s, w_out);
    input wire [31:0] w_in1, w_in2;
    input wire w_s;
    output wire [31:0] w_out;
    assign w_out = (w_s) ? w_in1 : w_in2;
endmodule