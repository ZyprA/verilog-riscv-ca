`default_nettype none

module m_am_imem(w_pc, w_inst);
    input wire [31:0] w_pc;
    output wire [31:0] w_inst;
    reg [31:0] mem [63:0];
    assign w_inst = mem[w_pc[7:2]];
    integer i; initial for (i=0; i<64; i=i+1) mem[i]=32'd0;
endmodule