`default_nettype none

module m_sm_dmem(w_clk, w_adr, w_we, w_wd, r_rd);
    input wire w_clk, w_we;
    input wire [31:0] w_adr, w_wd;
    output reg [31:0] r_rd;
    reg [31:0] mem [0:63];
    always @(posedge w_clk) r_rd <= mem[w_adr[7:2]];
    always @(posedge w_clk) if (w_we) mem[w_adr[7:2]] <= w_wd;
    integer i; initial for (i=0; i<64; i=i+1) mem[i] = 32'd0;
endmodule