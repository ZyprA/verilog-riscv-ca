`default_nettype none

module m_alu(w_in1, w_in2, w_out, w_tkn);
    input wire [31:0] w_in1, w_in2;
    output wire [31:0] w_out;
    output wire w_tkn;
    assign w_out = w_in1 + w_in2;
    assign w_tkn = (w_in1 != w_in2);
endmodule